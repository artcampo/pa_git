library ieee;
use ieee.std_logic_1164.all;
use work.proc_package.all;

package tb_load_signals is

signal p256           : std_logic_vector(data_width_c - 1 downto 0);	
signal p257           : std_logic_vector(data_width_c - 1 downto 0);	

end package tb_load_signals;