library ieee;
use ieee.std_logic_1164.all;
use work.proc_package.all;

package tb_load_signals is

signal p0           : std_logic_vector(data_width_c - 1 downto 0);	
signal p1           : std_logic_vector(data_width_c - 1 downto 0);	
signal p2           : std_logic_vector(data_width_c - 1 downto 0);	
signal p3           : std_logic_vector(data_width_c - 1 downto 0);	
signal p4           : std_logic_vector(data_width_c - 1 downto 0);	

end package tb_load_signals;