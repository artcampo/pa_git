library ieee;
use ieee.std_logic_1164.all;

package tb_package is

-------------------------------------------------------------------------------------



end package tb_package;